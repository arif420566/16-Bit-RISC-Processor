/*************************************************************
Design Name 	: 
File Name   	: .v
Function    	: 
Coder		    	: 
Last Modified	: 
*************************************************************/

module mux2_to_1(in0,in1,sel,out);
	input [15:0] in0,in1;
	input sel;
	output [15:0] out;

	reg [15:0] out;

	always @(sel or in0 or in1)
	begin
		case(sel)
			1'b0: out=in0;
			1'b1: out=in1;
		endcase
	end
	
endmodule
